`timescale 1ns/1ns
// Testbench for the VGA Module

module vga_tb();
//-- Setup parameters to pass to the DUT
localparam INTERFACE_WIDTH_BITS = 128;
localparam BITS_PER_PIXEL = 16;
localparam CLOCK_FREQ_HZ = 25_000_000;

//-- Should probably not change these.
localparam DISPLAY_WIDTH        = 640;
localparam DISPLAY_HEIGHT       = 480;
localparam INTERFACE_ADDR_BITS  = 26;

//-- Calculated parameters
// Use integer division here to avoid a pixel being split across two
// addresses in the buffer
localparam PIXELS_PER_TRANSFER = INTERFACE_WIDTH_BITS / BITS_PER_PIXEL;
localparam INTERFACE_WIDTH_BYTES = INTERFACE_WIDTH_BITS / 8;

// Use $ceil to ensure we get all pixels.
// Without $rtoi, NUM_BUFFER_ENTRIES ends up being a float which causes
// complications down the line as it is used to define the bit-widths of
// various signals.
localparam NUM_BUFFER_ENTRIES = $rtoi($ceil(DISPLAY_WIDTH / PIXELS_PER_TRANSFER));

//-- DUT Signals.
logic clk;
logic reset_n;

// VGA Timing Signals
logic [3:0] VGA_R, VGA_G, VGA_B;
logic VGA_HS, VGA_VS;

// Indicate display active.
logic display_enabled;

logic [INTERFACE_ADDR_BITS-1:0] image_base_address;
logic buffer_start;
logic [INTERFACE_ADDR_BITS-1:0]          buffer_base_address;
logic [$clog2(NUM_BUFFER_ENTRIES)-1:0]   buffer_read_addr;
logic [INTERFACE_WIDTH_BITS-1:0]          buffer_read_data;

logic end_frame;

// --------------- //
// Instantiate DUT //
// --------------- //
vga #(
    .INTERFACE_WIDTH_BITS   (INTERFACE_WIDTH_BITS),
    .BITS_PER_PIXEL         (BITS_PER_PIXEL),
    .DISPLAY_WIDTH          (DISPLAY_WIDTH),
    .DISPLAY_HEIGHT         (DISPLAY_HEIGHT),
    .NUM_BUFFER_ENTRIES     (NUM_BUFFER_ENTRIES),
    .INTERFACE_ADDR_BITS    (INTERFACE_ADDR_BITS)
) DUT (
    .clk        (clk),
    .reset_n    (reset_n),
    .VGA_R      (VGA_R),
    .VGA_G      (VGA_G),
    .VGA_B      (VGA_B),
    .VGA_HS     (VGA_HS),
    .VGA_VS     (VGA_VS),
    .display_enabled        (display_enabled),
    .image_base_address     (image_base_address),
    .buffer_start           (buffer_start),
    .buffer_base_address    (buffer_base_address),
    .buffer_read_addr       (buffer_read_addr),
    .buffer_read_data       (buffer_read_data),
    .end_frame              (end_frame)
);

//------------------------------------------------------------------------------
// The "ground-truth" pixel data will be stored in a global array in this test
// bench.
//
// Each time the VGA module generates a "start" signals, a buffer mimic will
// load data from this ground truth and service read requests from the DUT
// with a latency of one clock cycle.
//
// To verify the correctness of the module, the red, green, and blue signals
// will be concatenated together and compared against the lower 12 bits of the
// ground truth pixel buffer.

localparam NUM_PIXELS = DISPLAY_WIDTH * DISPLAY_HEIGHT;
logic [BITS_PER_PIXEL-1:0] pixels [NUM_PIXELS-1:0];

// Buffer mimic.
logic [INTERFACE_WIDTH_BITS-1:0] buffer [NUM_BUFFER_ENTRIES-1:0];

// -- Helper routines --

// Setup the clock
initial begin
    clk = 0;
    forever #(CLOCK_FREQ_HZ / 2) clk = ~clk;
end

// Turn a address reference generated by the DUT into an index into the
// "pixels" array.
//
// NOTE: image_base_address must be held constant throughout the entirety of
// a single frame.
function automatic int make_index;
    input [INTERFACE_ADDR_BITS-1:0] address;
    begin
        return (address - image_base_address) * PIXELS_PER_TRANSFER / INTERFACE_WIDTH_BYTES;
    end

endfunction


// Handle start requests by the DUT
always @(posedge buffer_start) begin : Load_Buffer
    automatic int index = make_index(buffer_base_address);
    //$display("index = %d", index);
    for (int i = 0; i < NUM_BUFFER_ENTRIES; i = i+1) begin
        for (int j = 0; j < PIXELS_PER_TRANSFER; j = j+1) begin
            // Pack pixel data into each entry in the buffer
            buffer[i][(BITS_PER_PIXEL * j) +: BITS_PER_PIXEL] = pixels[index];
            index = index + 1;
        end    
    end
end

// Handle read requests by the DUT
always @(posedge clk) begin
    buffer_read_data <= buffer[buffer_read_addr];
end

// Assign the reset signal.
task assert_reset();
    reset_n = 1'b0;
    @(posedge clk);
    reset_n = 1'b1;
endtask

// Main test loop
initial begin : Main_Test
    // Local signals
    logic [11:0] this_pixel;
    logic [11:0] expected_pixel;

    // Keep track of the number of cycles "display_enable" has been asserted
    // to track which pixel should be displayed. Used to check the validity of
    // the output.
    automatic int output_index;

    // Randomize the contents of the pixel data
    for (int i = 0; i < NUM_PIXELS; i = i+1) begin
        pixels[i] = $urandom();
    end 

    reset_n = 1'b1;
    image_base_address = 4'h1000;

    assert_reset();

    // Wait until the start of the first valid frame.
    @(posedge buffer_start);  
    @(posedge display_enabled);

    // Loop until all pixels should have been displayed.
    output_index = DISPLAY_WIDTH;
    while (output_index < NUM_PIXELS) begin
        // Wait until the negative edge of the clock. All signals should be
        // resolved by this point.
        @(negedge clk);
        
        if (display_enabled) begin
            this_pixel = {VGA_B, VGA_G, VGA_R};
            // Get the expected pixel from "pixels" array
            expected_pixel = pixels[output_index];
            assert(this_pixel == expected_pixel);

            // Prepare for the net pixel.
            output_index = output_index + 1; 
        end
    end

    // End simulation.
    $stop;
end


endmodule
